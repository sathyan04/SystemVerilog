module for_loop();
  int i;
  initial begin
    for(i=0;i<10;i++) begin
      $display("Iteration: %0d",i);
    end
  end
endmodule

/*
Output:

Iteration: 0
Iteration: 1
Iteration: 2
Iteration: 3
Iteration: 4
Iteration: 5
Iteration: 6
Iteration: 7
Iteration: 8
Iteration: 9

*/
